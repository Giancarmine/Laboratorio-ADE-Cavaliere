* C:\Users\hp\Documents\Laboratorio-ADE-Cavaliere\Latch SR\NOR Sync\NOR Sync.sch

* Schematics Version 9.1 - Web Update 1
* Wed May 06 15:44:55 2015



** Analysis setup **
.tran 0ns 1000ns


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "NOR Sync.net"
.INC "NOR Sync.als"


.probe


.END
