* C:\Users\hp\Documents\Laboratorio-ADE-Cavaliere\Latch SR\NOR Sync\NOR Sync.sch

* Schematics Version 9.1 - Web Update 1
* Thu May 07 10:57:32 2015



** Analysis setup **
.tran 0ns 1000ns


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "NOR Sync.net"
.INC "NOR Sync.als"


.probe


.END
