* C:\Users\hp\Documents\Laboratorio-ADE-Cavaliere\Latch SR\NAND Sync\NAND Sync.sch

* Schematics Version 9.1 - Web Update 1
* Thu May 07 12:15:03 2015



** Analysis setup **
.tran 0ns 1000ns


* From [PSPICE NETLIST] section of pspiceev.ini:
.lib "nom.lib"

.INC "NAND Sync.net"
.INC "NAND Sync.als"


.probe


.END
